library ieee;use ieee.std_logic_1164.all;use ieee.std_logic_unsigned.all;entity Johnson_counter is	port (		clk: in std_logic;		data_out: out std_logic_vector(3 downto 0)	);end Johnson_counter;architecture Johnson_counter_part of Johnson_counter issignal drop: std_logic_vector(3 downto 0);signal data_list: std_logic_vector(4 downto 0);component Johnson_D is	port (		clk, d: in std_logic;		q: inout std_logic;		not_q: out std_logic	);end component;begin	data_list(0) <= drop(3);	forloop1: for i in 0 to 3 generate		Johnson: Johnson_D port map(clk, data_list(i), data_list(i+1), drop(i));		data_out(i) <= data_list(i+1);	end generate forloop1;end Johnson_counter_part;